`ifndef TVIP_AXI_STATUS_SVH
`define TVIP_AXI_STATUS_SVH
class tvip_axi_status extends tue_status;
  `tue_object_default_constructor(tvip_axi_status)
  `uvm_object_utils(tvip_axi_status)
endclass
`endif
