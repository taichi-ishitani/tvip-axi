`ifndef TVIP_AXI_MASTER_RAL_PREDICTOR_SVH
`define TVIP_AXI_MASTER_RAL_PREDICTOR_SVH
typedef uvm_reg_predictor #(tvip_axi_master_item) tvip_axi_master_ral_predictor;
`endif
